library verilog;
use verilog.vl_types.all;
entity inccomp2 is
end inccomp2;
