module instr_mem (
	clk,
	memRead,
	memWrite,
	address,
	imem_in,
	imem_out
	);

input  clk, memRead, memWrite;
input [6:0] address;
input [31:0] imem_in;
output [31:0] imem_out;

reg [31:0] imem_out;

always @ (posedge clk)
begin
	imem_out = 32'b00000000000000000000000000000000;
	if (memRead) begin
		case (address)
			7'b0000000 : imem_out = 32'b00000000011100000000100000010011;
			7'b0000100 : imem_out = 32'b00000000000000000010001000010111;
			7'b0001000 : imem_out = 32'b11111111110000100000001000010011;
			7'b0001100 : imem_out = 32'b00000000000000000010001010010111;
			7'b0010000 : imem_out = 32'b00000001000000101000001010010011;
			7'b0010100 : imem_out = 32'b01000000000000000000011010110111;
			7'b0011000 : imem_out = 32'b11111111111101101000011010010011;
			7'b0011100 : imem_out = 32'b00000010000010000000100001100011;
			7'b0100000 : imem_out = 32'b00000000000000100010010000000011;
			7'b0100100 : imem_out = 32'b01000001111101000101010010010011;
			7'b0101000 : imem_out = 32'b00000000100101000100010100110011;
			7'b0101100 : imem_out = 32'b00000000000101001111010010010011;
			7'b0110000 : imem_out = 32'b00000000100101010000010100110011;
			7'b0110100 : imem_out = 32'b00000000010000100000001000010011;
			7'b0111000 : imem_out = 32'b11111111111110000000100000010011;
			7'b0111100 : imem_out = 32'b00000000110101010010010110110011;
			7'b1000000 : imem_out = 32'b11111100000001011000111011100011;
			7'b1000100 : imem_out = 32'b00000000000001010000011010110011;
			7'b1001000 : imem_out = 32'b11111101010111111111000011101111;
			7'b1001100 : imem_out = 32'b00000000110100101010000000100011;
			7'b1010000 : imem_out = 32'b00000000000000000000000011101111;
			7'b1010100 : imem_out = 32'b00000000000000000000000000010011;
		endcase
	end
end

endmodule